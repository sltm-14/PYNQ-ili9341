`ifndef pkg_loop
`define pkg_loop

package pkg_loop;



endpackage
`endif
