library verilog;
use verilog.vl_types.all;
entity pkg_ili9341 is
end pkg_ili9341;
