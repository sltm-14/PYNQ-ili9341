library verilog;
use verilog.vl_types.all;
entity pkg_loop is
end pkg_loop;
