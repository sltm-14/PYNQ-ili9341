library verilog;
use verilog.vl_types.all;
entity send_command_sv_unit is
end send_command_sv_unit;
